library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity robot is
    port (
        clk             : in std_logic;
        reset           : in std_logic;
        
        sensor_l_in     : in std_logic;  
        sensor_m_in     : in std_logic;       
        sensor_r_in     : in std_logic;

        motor_l_pwm     : out std_logic;
        motor_r_pwm     : out std_logic;       
        
        mine_square_in  : in std_logic;
        ro_rx              : in std_logic; 
        ro_tx              : out std_logic;

        treasure_sw         : in std_logic;
		  
		  DEB_led : out std_logic_vector(6 downto 0)
    );
end entity robot;

architecture structural of robot is
    component controller is
        port (
            sensors_out	        : in std_logic_vector (2 downto 0); 
            clk	                : in std_logic;
            reset	   	        : in std_logic;
            count_in    	    : in std_logic_vector (19 downto 0);
            ctr_mine            : in std_logic;
            ctr_data            : in std_logic_vector (7 downto 0);

            int_count_ctrl      : in std_logic_vector (31 downto 0);
            int_reset_ctrl      : out std_logic;

            treasure_sw         : in std_logic;
            
            count_reset         : out std_logic;
            direction_l	        : out std_logic;	
            direction_l_reset   : out std_logic;
            direction_r         : out std_logic;
            direction_r_reset   : out std_logic;
            ctr_mine_out        : out std_logic;
            ctr_mid             : out std_logic;
				
				DEB_led : out std_logic_vector(4 downto 0);
				  led_DEB :out std_logic_vector(1 downto 0)
    
      );
    end component controller;

    component eightbitregister is
        port(             
            clk                     :in std_logic;  
				reset							:in std_logic;
            register_input          :in std_logic_vector(7 downto 0);
    
            register_output         :out std_logic_vector(7 downto 0)
    );
    end component eightbitregister;

    component Data_sender is
        port (
            clk             : in std_logic;
            reset           : in std_logic;
        -- tx
            DS_out_UART_in  : out std_logic_vector(7 downto 0);
            buffer_empty    : in std_logic;
            DS_write           : out std_logic;
        -- rx
            DS_in_UART_out  : in std_logic_vector(7 downto 0);
            data_ready      : in std_logic;
            DS_read            : out std_logic;
        -- user in
            DS_in_mine      : in std_logic;
            DS_in_mid       : in std_logic;
            DS_out          : out std_logic_vector(7 downto 0)
      );
    end component Data_sender;

    component Mine_detector is
        generic (
            trig_count      : integer := 2700 -- (50*10^6/trig_freq)/2
            );
          port (
            clk             : in std_logic;
            reset           : in std_logic;
            square_in       : in std_logic;
            sensors_out     : in std_logic_vector(2 downto 0);
            register_output : in std_logic_vector (8 downto 0);
            
            mine_out        : out std_logic;
            register_input : out std_logic_vector(8 downto 0);
            register_enable : out std_logic
          );
    end component Mine_detector;

    component eightbitmemory is
        port(   register_input       :in std_logic_vector(8 downto 0);
                clk         :in std_logic;
                reset			: in std_logic;
    
                enable	: in std_logic;
                register_output      :out std_logic_vector(8 downto 0)
        );
    end component eightbitmemory;

    component motorcontrol is
        port (
        reset			: in	std_logic;
        direction		: in	std_logic;
        count_in		: in	std_logic_vector (19 downto 0);
        pwm			    : out	std_logic :='1'
        );
    end component motorcontrol;

    component inputbuffer is
        port(
            clk                 : in std_logic;
            sensor_l_in         : in std_logic;
            sensor_m_in         : in std_logic; 
            sensor_r_in         : in std_logic;
            sensors_out         : out std_logic_vector(2 downto 0)
        );
    end component inputbuffer;

    component timebase is
        port(
            clk                     : in std_logic;
            reset                   : in std_logic;
            count_out               : out std_logic_vector(19 downto 0)
        );
    end component timebase;

    component IntegerOfTime is
        port (clk                   : in std_logic;
              reset                 : in std_logic;
              int_count_out         : out std_logic_vector(31 downto 0)
        );
        end component IntegerOfTime;

    component uart is
        port (
            clk             : in  std_logic;
            reset           : in  std_logic;
    
            rx              : in  std_logic;
            tx              : out std_logic;
    
            data_in         : in  std_logic_vector (7 downto 0);
            buffer_empty    : out std_logic;
            write           : in  std_logic;
    
            data_out        : out std_logic_vector (7 downto 0);
            data_ready      : out std_logic;
            read            : in  std_logic
        );
    end component uart;

    signal direction_ll, direction_l_resett, direction_rr, direction_r_resett       : std_logic;
    signal count                                                                    : std_logic_vector (19 downto 0);
    signal int_count                                                                : std_logic_vector (31 downto 0);
    signal reset_counter, Int_Count_reset                                           : std_logic;                         
    --Internal reset for counter and such
    signal sensors_out                                                              : std_logic_vector (2 downto 0);
    signal mine_detect_ctr, mine_detect_ds                                          : std_logic; 
    signal data_in, data_out                                                        : std_logic_vector (7 downto 0); 
    signal ds_in_mid_s, read_s, data_ready_s, buffer_empty_s, write_s               : std_logic;
    signal ds_out_uart_in_s, DS_in_UART_out_s                                       : std_logic_vector (7 downto 0);
    signal mine_mem_in_sig, mine_mem_out_s                                          : std_logic_vector (8 downto 0);
    signal mem_en                                                                   : std_logic; 
begin
    -- external signal handling

    CRT: controller port map(
                                sensors_out     	=> sensors_out,                           
                                clk     		    => clk,
                                reset             	=> reset,
                                count_in     		=> count,
                                ctr_mine            => mine_detect_ctr,
                                ctr_data            => data_out,

                                int_count_ctrl => int_count,
                                int_reset_ctrl => Int_Count_reset,

                                treasure_sw => treasure_sw,

                                count_reset     	=> reset_counter,
                                direction_l     	=> direction_ll,
                                direction_l_reset   => direction_l_resett,
                                direction_r     	=> direction_rr,
                                direction_r_reset   => direction_r_resett,
                                ctr_mine_out        => mine_detect_ds,
                                ctr_mid             => ds_in_mid_s,
										  
										  DEB_led(0) => DEB_led(0),
										  DEB_led(1) => DEB_led(1),
										  DEB_led(2) => DEB_led(2),
										  DEB_led(3) => DEB_led(3),
										  DEB_led(4) => DEB_led(4),
										  led_DEB(0) => DEB_led(5),
										  led_DEB(1) =>DEB_led(6)
										  
    );

    REG: eightbitregister port map(
                                clk                 => clk,
										  reset					 => reset,
                                register_input      => data_in,

                                register_output     => data_out
    );

    DS: data_sender port map(      
                                clk                 => clk,
                                reset               => reset,
                            -- tx          =>
                                DS_out_UART_in      =>  ds_out_uart_in_s,
                                buffer_empty        =>  buffer_empty_s,
                                DS_write               =>  write_s,
                            -- rx      =>
                                DS_in_UART_out      =>  DS_in_UART_out_s,   
                                data_ready          =>  data_ready_s,
                                DS_read                =>  read_s,
                            -- user in     =>
                                DS_in_mine          =>  mine_detect_ds,
                                DS_in_mid           =>  ds_in_mid_s,
                                DS_out              =>  data_in
                            
    );    

    MD: Mine_detector port map (
                                clk                => clk,
                                reset              => reset,
                                square_in          => mine_square_in,
                                sensors_out        => sensors_out,
                                register_output    <= mine_mem_out_s,

                                mine_out           => mine_detect_ctr,
                                register_input     => mine_mem_in_sig,
                                register_enable    => mine_mem_out_s

    MEM: eightbitmemory port map (
                                register_input      <= mine_mem_in_sig,
                                clk                 => clk,
                                reset			    => reset,

                                enable	            <= mem_en,
                                register_output     => mine_mem_out_s
    );

    MCL: motorcontrol port map(
                                reset               => direction_l_resett,
                                direction           => direction_ll,
                                count_in            => count,

                                pwm                 => motor_l_pwm
    );

    MCR: motorcontrol port map(
                                reset               => direction_r_resett,
                                direction           => direction_rr,
                                count_in            => count,

                                pwm                 => motor_r_pwm
    );

    IB: inputbuffer port map(
                                clk                 => clk,
                                sensor_l_in         => sensor_l_in,
                                sensor_m_in         => sensor_m_in,
                                sensor_r_in         => sensor_r_in,

                                sensors_out         => sensors_out
    );

    TB: timebase port map(
                                clk                 => clk,
                                reset               => reset_counter,

                                count_out           => count
    );

    ITB: IntegerOfTime port map (
                  clk                   => clk,
                  reset                 => Int_Count_reset,
                  int_count_out         => int_count
    );

    ua : UART port map(
                                clk                 => clk,
                                reset               => reset,

                                rx                  =>  ro_rx,
                                tx                  =>  ro_tx,

                                data_in             => ds_out_uart_in_s,
                                buffer_empty        => buffer_empty_s,
                                write               => write_s,

                                data_out            => DS_in_UART_out_s,
                                data_ready          => data_ready_s,
                                read                => read_s
    );
    
    
end architecture structural;
